module UartTxrTB();

endmodule
